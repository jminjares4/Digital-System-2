`timescale 1ns / 1ps

module Lab3tb;

endmodule
